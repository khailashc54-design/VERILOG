module srlatch(input s,r, output q,qbar);
  assign q=~(~r&qbar);
  assign qbar=~(~s&q);
endmodule


module srlatch_tb;
  reg s,r;
  wire q,qbar;
  srlatch dut(.*);
  initial begin
  $monitor("t=%0t|s=%b r=%b|q=%b qbar=%b",$time,s,r,q,qbar);
  s=0;r=0;
  #10 s=1;r=0;
  #10 s=0;r=1;
  #10 s=1;r=1;
  $finish;
  end
  endmodule

